library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity template is
	port (
		clk : in std_logic;
		rst : in std_logic;
		sig
	);
end template;

architecture rtl of template is

begin

end architecture;